module data

fn test_max() {
    arr := [3, 5, 1, 2 ]
    high := max(arr)
    assert high == 5
}

